.title KiCad schematic
C1 Net-_C1-Pad1_ 0 1u
C2 out 0 100n
V1 Net-_V1-E1_ 0 dc 0 pulse (0 5 1u 1u 1u 1 1)
R2 Net-_C1-Pad1_ out 1k
R1 Net-_V1-E1_ Net-_C1-Pad1_ 10k
.tran 50u 50m
.end

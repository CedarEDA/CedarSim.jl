*My Title
.GLOBAL VDD
.GLOBAL VSS
VVDD VDD 0 5.0
VVSS VSS 0 0.0
.END

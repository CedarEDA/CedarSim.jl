.param gmin=1e-15
.OPTION afsmode=5 parasitics=1
.OPT gmin=gmin donominal=1
.OPTIONS montecon=1 montemeas=1 montequantiles=[0.134989803163 99.865010196837]
.OPTIONS REMOVEVSRC=0 STATFL=1
.OPT LISLVL=1 NOMOD SYMB=1 POST_VERSION=2001
.OPTION POST PROBE
.OPTIONS NUMDGT=10 MEASDGT=10 AUTOSTOP OPTS
.width out = 256
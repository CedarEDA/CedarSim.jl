m0 d1 g s1 b nmos_3p3 W=1e-6 l=1e-6

 .param
 +nmos_3p3_noia='3.2e+041 + 3.5e+042' 
 +nmos_3p3_noib='1.2e+020 + 1.2e+020' 
 +nmos_3p3_noic='6.0e+008 + 6.0e+008'
.model  nmos_3p3.0  nmos
+level = 54
+lmin    = 2.8e-007      
+lmax    = 5e-007        
+wmin    = 2.2e-007      
+wmax    = 5e-007        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.70837662    
+lvth0   = -3.8715455e-008
+wvth0   = -1.430587e-008
+pvth0   = 4.3636364e-016
+k1      = 0.95938091    
+lk1     = -9.9985454e-008
+k2      = 0.054714558   
+lk2     = -4.1647636e-008
+wk2     = -1.9242857e-008
+pk2     = 5.388e-015    
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.1262652    
+lvoff   = 3.9354545e-009
+wvoff   = 5.3064935e-009
+pvoff   = -1.4858182e-015
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.023671338   
+lu0     = 4.6525455e-009
+wu0     = 4.6066597e-009
+pu0     = -6.5127273e-016
+ua      = -1.1554452e-009
+lua     = 7.0220545e-016
+wua     = 2.7073777e-016
+pua     = -1.4149745e-022
+ub      = 3.3771156e-018
+lub     = -7.9058636e-025
+wub     = -4.093733e-025
+pub     = 9.2644364e-032
+uc      = 2.2660166e-010
+luc     = -6.1360545e-017
+wuc     = -3.2577351e-017
+puc     = 5.4467782e-024
+eu      = 1.67          
+vsat    = 92454.546     
+lvsat   = -0.0027272727 
+wvsat   = -0.00021818182
+pvsat   = 1.3090909e-009
+a0      = 0.11197377    
+la0     = -3.1454545e-009
+wa0     = -6.2322078e-009
+pa0     = 1.7450182e-015
+ags     = 0.32403844    
+lags    = -1.5116364e-008
+wags    = 4.7930493e-008
+pags    = -1.2213818e-014
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.14896036   
+lketa   = 3.8830182e-008
+wketa   = 8.1643636e-009
+pketa   = -2.4261818e-015
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.3741        
+lpclm   = -4.729e-008   
+wpclm   = 2.1028364e-008
+ppclm   = 8.5658182e-015
+pdiblc1 = 0.39          
+pdiblc2 = 0.003171      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0036363636  
+ldelta  = 3.1818182e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 2.652013e-006 
+lalpha0 = -3.0506364e-013
+walpha0 = 4.8779221e-014
+palpha0 = -1.3658182e-020
+alpha1  = 0             
+beta0   = 19.905584     
+lbeta0  = 1.2863636e-007
+wbeta0  = 1.3848312e-007
+pbeta0  = 8.7272727e-016
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.45934558   
+lkt1    = 4.2126364e-008
+wkt1    = 3.2086753e-008
+pkt1    = -8.6530909e-015
+kt1l    = 0             
+kt2     = -0.024730519  
+lkt2    = 1.2545455e-009
+wkt2    = 1.0597403e-009
+pkt2    = -2.9672727e-016
+ute     = -1.5675325    
+lute    = 9.0909091e-008
+wute    = 1.0441558e-007
+pute    = -4.3636364e-014
+ua1     = 1.675e-009    
+ub1     = -4.1945234e-018
+lub1    = 2.8745455e-025
+wub1    = 3.3492467e-025
+pub1    = -5.7490909e-032
+uc1     = -4.2363636e-011
+luc1    = -3.8181818e-018
+wuc1    = -6.5454545e-018
+puc1    = 1.8327273e-024
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.1  nmos
+level = 54
+lmin    = 5e-007        
+lmax    = 1.2e-006      
+wmin    = 2.2e-007      
+wmax    = 5e-007        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.67781184    
+lvth0   = -2.3433061e-008
+wvth0   = -1.2304653e-008
+pvth0   = -5.642449e-016
+k1      = 0.74639857    
+lk1     = 6.5057143e-009
+k2      = 0.0237458     
+lk2     = -2.6163257e-008
+wk2     = -3.01296e-009 
+pk2     = -2.7269486e-015
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.11273959   
+lvoff   = -2.8273469e-009
+wvoff   = 1.6942041e-009
+pvoff   = 3.2032653e-016
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.029675694   
+lu0     = 1.6503673e-009
+wu0     = 8.572898e-010 
+pu0     = 1.2234122e-015
+ua      = -1.2961984e-009
+lua     = 7.7258204e-016
+wua     = 4.7264816e-017
+pua     = -2.976098e-023
+ub      = 3.0836898e-018
+lub     = -6.4387347e-025
+wub     = -2.7080816e-026
+pub     = -9.8501878e-032
+uc      = 8.4613959e-011
+luc     = 9.6333061e-018
+wuc     = 2.2398367e-018
+puc     = -1.1961815e-023
+eu      = 1.67          
+vsat    = 83571.429     
+lvsat   = 0.0017142857  
+wvsat   = -0.0017142857 
+pvsat   = 2.0571429e-009
+a0      = 1.0861147     
+la0     = -4.9021592e-007
+wa0     = -5.1997224e-008
+pa0     = 2.4627526e-014
+ags     = 0.47870122    
+lags    = -9.2447755e-008
+wags    = 4.3304327e-008
+pags    = -9.9007347e-015
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.028417143  
+lketa   = -2.1441429e-008
+wketa   = -7.4262857e-009
+pketa   = 5.3691429e-015
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.082893878   
+lpclm   = 9.8313061e-008
+wpclm   = 4.3902367e-008
+ppclm   = -2.8711837e-015
+pdiblc1 = 0.39          
+pdiblc2 = 0.001359      
+lpdiblc2= 9.06e-010     
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0014285714  
+ldelta  = 4.2857143e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 6.5720816e-006
+lalpha0 = -2.265098e-012
+walpha0 = -1.5330612e-014
+palpha0 = 1.8396735e-020
+alpha1  = 0             
+beta0   = 22.625306     
+lbeta0  = -1.2312245e-006
+wbeta0  = -3.5054694e-007
+pbeta0  = 2.4538775e-013
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.33916633   
+lkt1    = -1.7963265e-008
+wkt1    = -2.4641633e-009
+pkt1    = 8.6223674e-015
+kt1l    = 0             
+kt2     = -0.020311225  
+lkt2    = -9.5510204e-010
+wkt2    = -3.9183673e-011
+pkt2    = 2.5273469e-016
+ute     = -1.3857143    
+wute    = 1.7142857e-008
+ua1     = 1.675e-009    
+ub1     = -2.804398e-018
+lub1    = -4.0760816e-025
+wub1    = 5.6899592e-026
+pub1    = 8.1521633e-032
+uc1     = -6.0285714e-011
+luc1    = 5.1428571e-018
+wuc1    = 2.0571429e-018
+puc1    = -2.4685714e-024
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.2  nmos
+level = 54
+lmin    = 1.2e-006      
+lmax    = 1e-005        
+wmin    = 2.2e-007      
+wmax    = 5e-007        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.66097097    
+lvth0   = -3.224026e-009
+wvth0   = -9.7008312e-009
+pvth0   = -3.6888312e-015
+k1      = 0.79593364    
+lk1     = -5.2936364e-008
+k2      = 0.0056393844  
+lk2     = -4.4355584e-009
+wk2     = -7.4596769e-009
+pk2     = 2.6091117e-015
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12631325   
+lvoff   = 1.3461039e-008
+wvoff   = 2.0819221e-009
+pvoff   = -1.4493507e-016
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.032447266   
+lu0     = -1.6755195e-009
+wu0     = 6.7095584e-010
+pu0     = 1.447013e-015 
+ua      = -8.1547091e-010
+lua     = 1.9570909e-016
+wua     = 6.0458182e-018
+pua     = 1.9701818e-023
+ub      = 2.7427942e-018
+lub     = -2.347987e-025
+wub     = -1.6048831e-026
+pub     = -1.1174026e-031
+uc      = 9.84685e-011  
+luc     = -6.9921429e-018
+wuc     = -8.8975636e-018
+puc     = 1.4030649e-024
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.224418      
+la0     = -6.5617987e-007
+wa0     = 4.291948e-009 
+pa0     = -4.2919481e-014
+ags     = 0.25784649    
+lags    = 1.7257792e-007
+wags    = -2.606026e-009
+pags    = 4.5191688e-014
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.019651071  
+lketa   = -3.1960714e-008
+wketa   = -6.5992208e-010
+pketa   = -2.7504935e-015
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.18918506    
+lpclm   = -2.9236364e-008
+wpclm   = 2.1551688e-009
+ppclm   = 4.7225454e-014
+pdiblc1 = 0.39          
+pdiblc2 = 0.00064013636 
+lpdiblc2= 1.7686364e-009
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0027272727  
+ldelta  = 2.7272727e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 7.5243347e-005
+lalpha0 = -8.4670617e-011
+walpha0 = 7.5358442e-012
+palpha0 = -9.043013e-018
+alpha1  = 0             
+beta0   = 24.210162     
+lbeta0  = -3.133052e-006
+wbeta0  = 1.1381299e-007
+pbeta0  = -3.1184416e-013
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.32898149   
+lkt1    = -3.0185065e-008
+wkt1    = -7.3528831e-009
+pkt1    = 1.4488831e-014
+kt1l    = 0             
+kt2     = -0.021107143  
+wkt2    = 1.7142857e-010
+ute     = -1.3857143    
+wute    = 1.7142857e-008
+ua1     = 1.675e-009    
+ub1     = -2.5166039e-018
+lub1    = -7.5296104e-025
+wub1    = 2.224987e-026 
+pub1    = 1.231013e-031 
+uc1     = -5.6e-011     
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.3  nmos
+level = 54
+lmin    = 1e-005        
+lmax    = 5.0001e-005   
+wmin    = 2.2e-007      
+wmax    = 5e-007        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.66064857    
+wvth0   = -1.0069714e-008
+k1      = 0.79064       
+k2      = 0.0051958286  
+wk2     = -7.1987657e-009
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12496714   
+wvoff   = 2.0674286e-009
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.032279714   
+wu0     = 8.1565714e-010
+ua      = -7.959e-010   
+wua     = 8.016e-018    
+ub      = 2.7193143e-018
+wub     = -2.7222857e-026
+uc      = 9.7769286e-011
+wuc     = -8.7572571e-018
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.1588        
+ags     = 0.27510429    
+wags    = 1.9131429e-009
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.022847143  
+wketa   = -9.3497143e-010
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.18626143    
+wpclm   = 6.8777143e-009
+pdiblc1 = 0.39          
+pdiblc2 = 0.000817      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.003         
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 6.6776286e-005
+walpha0 = 6.6315429e-012
+alpha1  = 0             
+beta0   = 23.896857     
+wbeta0  = 8.2628571e-008
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.332        
+wkt1    = -5.904e-009   
+kt1l    = 0             
+kt2     = -0.021107143  
+wkt2    = 1.7142857e-010
+ute     = -1.3857143    
+wute    = 1.7142857e-008
+ua1     = 1.675e-009    
+ub1     = -2.5919e-018  
+wub1    = 3.456e-026    
+uc1     = -5.6e-011     
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.4  nmos
+level = 54
+lmin    = 2.8e-007      
+lmax    = 5e-007        
+wmin    = 5e-007        
+wmax    = 1.2e-006      
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.72356597    
+lvth0   = -4.1979273e-008
+wvth0   = -2.1596758e-008
+pvth0   = 2.0029964e-015
+k1      = 0.95938091    
+lk1     = -9.9985454e-008
+k2      = 0.041255727   
+lk2     = -3.7879164e-008
+wk2     = -1.2782618e-008
+pk2     = 3.5791331e-015
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.079311948  
+lvoff   = -9.2114546e-009
+wvoff   = -1.7231065e-008
+pvoff   = 4.8246982e-015
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.033011551   
+lu0     = 4.0251818e-009
+wu0     = 1.2335751e-010
+pu0     = -3.5013818e-016
+ua      = -6.3005701e-010
+lua     = 3.9938436e-016
+wua     = 1.8551439e-017
+pua     = 3.8566691e-024
+ub      = 2.2836418e-018
+lub     = -9.0230909e-026
+wub     = 1.1549411e-025
+pub     = -2.4352626e-031
+uc      = 1.5877203e-010
+luc     = -3.4349127e-017
+wuc     = -1.9125195e-020
+puc     = -7.5187026e-024
+eu      = 1.67          
+vsat    = 71618.182     
+lvsat   = 0.0042909091  
+wvsat   = 0.0097832727  
+pvsat   = -2.0596364e-009
+a0      = 0.10680558    
+la0     = -1.6983636e-009
+wa0     = -3.7514805e-009
+pa0     = 1.0504145e-015
+ags     = 0.35500309    
+lags    = -1.1780546e-008
+wags    = 3.3067462e-008
+pags    = -1.3815011e-014
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.12490989   
+lketa   = 3.0254945e-008
+wketa   = -3.3798633e-009
+pketa   = 1.6899316e-015
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.45921829    
+lpclm   = -8.0088e-008  
+wpclm   = -1.9828414e-008
+ppclm   = 2.4308858e-014
+pdiblc1 = 0.39          
+pdiblc2 = 0.003171      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0036363636  
+ldelta  = 3.1818182e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 2.6500109e-006
+lalpha0 = -2.8170545e-013
+walpha0 = 4.9740218e-014
+palpha0 = -2.4870109e-020
+alpha1  = 0             
+beta0   = 20.982852     
+lbeta0  = -8.9454546e-008
+wbeta0  = -3.786053e-007
+pbeta0  = 1.0555636e-013
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.37773746   
+lkt1    = 1.6718727e-008
+wkt1    = -7.0851491e-009
+pkt1    = 3.5425745e-015
+kt1l    = 0             
+kt2     = -0.014603854  
+lkt2    = -3.3230727e-009
+wkt2    = -3.8010589e-009
+pkt2    = 1.9005294e-015
+ute     = -1.4342857    
+wute    = 4.0457143e-008
+ua1     = 1.675e-009    
+ub1     = -3.65896e-018 
+lub1    = 2.4878e-025   
+wub1    = 7.7854254e-026
+pub1    = -3.8927127e-032
+uc1     = -5.6e-011     
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.5  nmos
+level = 54
+lmin    = 5e-007        
+lmax    = 1.2e-006      
+wmin    = 5e-007        
+wmax    = 1.2e-006      
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.67504024    
+lvth0   = -1.7716408e-008
+wvth0   = -1.0974289e-008
+pvth0   = -3.3082384e-015
+k1      = 0.76833212    
+lk1     = -4.4610612e-009
+wk1     = -1.0528104e-008
+pk1     = 5.2640522e-015
+k2      = 0.0082103273  
+lk2     = -2.1356464e-008
+wk2     = 4.4440669e-009
+pk2     = -5.0342094e-015
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12049225   
+lvoff   = 1.1378694e-008
+wvoff   = 5.4154776e-009
+pvoff   = -6.4985731e-015
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.031181163   
+lu0     = 4.9403755e-009
+wu0     = 1.3466449e-010
+pu0     = -3.5579167e-016
+ua      = -1.1586455e-009
+lua     = 6.6367861e-016
+wua     = -1.8760555e-017
+pua     = 2.2512666e-023
+ub      = 2.8240225e-018
+lub     = -3.6042122e-025
+wub     = 9.755951e-026 
+pub     = -2.3455895e-031
+uc      = 8.1997037e-011
+luc     = 4.0383673e-018
+wuc     = 3.4959595e-018
+puc     = -9.2762449e-024
+eu      = 1.67          
+vsat    = 88428.571     
+lvsat   = -0.0041142857 
+wvsat   = -0.0040457143 
+pvsat   = 4.8548571e-009
+a0      = 0.97533082    
+la0     = -4.3596098e-007
+wa0     = 1.1790367e-009
+pa0     = -1.4148441e-015
+ags     = 0.441074      
+lags    = -5.4816e-008  
+wags    = 6.1365394e-008
+pags    = -2.7963977e-014
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.043888571  
+lketa   = -1.0255714e-008
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.21719837    
+lpclm   = 4.0921959e-008
+wpclm   = -2.0563788e-008
+ppclm   = 2.4676545e-014
+pdiblc1 = 0.39          
+pdiblc2 = 0.001359      
+lpdiblc2= 9.06e-010     
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0014285714  
+ldelta  = 4.2857143e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 6.8164074e-006
+lalpha0 = -2.3649037e-012
+walpha0 = -1.3260696e-013
+palpha0 = 6.6303478e-020
+alpha1  = 0             
+beta0   = 21.036008     
+lbeta0  = -1.1603265e-007
+wbeta0  = 4.1231608e-007
+pbeta0  = -2.8990433e-013
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.4079911    
+lkt1    = 3.1845551e-008
+wkt1    = 3.0571729e-008
+pkt1    = -1.5285865e-014
+kt1l    = 0             
+kt2     = -0.031229592  
+lkt2    = 4.9897959e-009
+wkt2    = 5.2016327e-009
+pkt2    = -2.6008163e-015
+ute     = -1.4342857    
+wute    = 4.0457143e-008
+ua1     = 1.675e-009    
+ub1     = -2.8098294e-018
+lub1    = -1.7578531e-025
+wub1    = 5.9506678e-026
+pub1    = -2.9753339e-032
+uc1     = -1.1888774e-010
+luc1    = 3.1443869e-017
+wuc1    = 3.0186115e-017
+puc1    = -1.5093057e-023
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.6  nmos
+level = 54
+lmin    = 1.2e-006      
+lmax    = 1e-005        
+wmin    = 5e-007        
+wmax    = 1.2e-006      
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.64923469    
+lvth0   = 1.325026e-008 
+wvth0   = -4.067414e-009
+pvth0   = -1.1596488e-014
+k1      = 0.79418892    
+lk1     = -3.5489221e-008
+wk1     = 8.3746286e-010
+pk1     = -8.3746286e-015
+k2      = -0.0057236965 
+lk2     = -4.6356351e-009
+wk2     = -2.005398e-009
+pk2     = 2.7051485e-015
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12197591   
+lvoff   = 1.3159091e-008
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.036490513   
+lu0     = -1.4308442e-009
+wu0     = -1.2698026e-009
+pu0     = 1.3295688e-015
+ua      = -7.881063e-010
+lua     = 2.1903156e-016
+wua     = -7.0891948e-018
+pua     = 8.5070338e-024
+ub      = 3.0594896e-018
+lub     = -6.4298182e-025
+wub     = -1.6806265e-025
+pub     = 8.4187636e-032
+uc      = 9.7557278e-011
+luc     = -1.4633922e-017
+wuc     = -8.460177e-018
+puc     = 5.071119e-024 
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.2333595     
+la0     = -7.4559545e-007
+ags     = 0.28370796    
+lags    = 1.3402325e-007
+wags    = -1.501953e-008
+pags    = 6.3697932e-014
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.021025909  
+lketa   = -3.7690909e-008
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.22708279    
+lpclm   = 2.9060649e-008
+wpclm   = -1.603574e-008
+ppclm   = 1.9242888e-014
+pdiblc1 = 0.39          
+pdiblc2 = 0.00064013636 
+lpdiblc2= 1.7686364e-009
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0027272727  
+ldelta  = 2.7272727e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 9.0921047e-005
+lalpha0 = -1.0329047e-010
+walpha0 = 1.0548281e-014
+palpha0 = -1.0548281e-019
+alpha1  = 0             
+beta0   = 24.039866     
+lbeta0  = -3.7206623e-006
+wbeta0  = 1.9555512e-007
+pbeta0  = -2.9791169e-014
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.33923366   
+lkt1    = -5.0663377e-008
+wkt1    = -2.4318421e-009
+pkt1    = 2.4318421e-014
+kt1l    = 0             
+kt2     = -0.021803571  
+lkt2    = -6.3214286e-009
+wkt2    = 5.0571429e-010
+pkt2    = 3.0342857e-015
+ute     = -1.7216234    
+lute    = 3.448052e-007 
+wute    = 1.7837922e-007
+pute    = -1.6550649e-013
+ua1     = 1.675e-009    
+ub1     = -3.5465249e-018
+lub1    = 7.0824935e-025
+wub1    = 5.1661197e-025
+pub1    = -5.7827969e-031
+uc1     = -5.0997566e-011
+luc1    = -5.0024338e-017
+wuc1    = -2.4011682e-018
+puc1    = 2.4011682e-023
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.7  nmos
+level = 54
+lmin    = 1e-005        
+lmax    = 5.0001e-005   
+wmin    = 5e-007        
+wmax    = 1.2e-006      
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.65055971    
+wvth0   = -5.2270629e-009
+k1      = 0.79064       
+k2      = -0.00618726   
+wk2     = -1.7348832e-009
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12066      
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.036347429   
+wu0     = -1.1368457e-009
+ua      = -7.6620314e-010
+wua     = -6.2384914e-018
+ub      = 2.9951914e-018
+wub     = -1.5964389e-025
+uc      = 9.6093886e-011
+wuc     = -7.9530651e-018
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.1588        
+ags     = 0.29711029    
+wags    = -8.6497371e-009
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.024795     
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.22998886    
+wpclm   = -1.4111451e-008
+pdiblc1 = 0.39          
+pdiblc2 = 0.000817      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.003         
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 8.0592e-005   
+alpha1  = 0             
+beta0   = 23.6678       
+wbeta0  = 1.92576e-007  
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.3443       
+kt1l    = 0             
+kt2     = -0.022435714  
+wkt2    = 8.0914286e-010
+ute     = -1.6871429    
+wute    = 1.6182857e-007
+ua1     = 1.675e-009    
+ub1     = -3.4757e-018  
+wub1    = 4.58784e-025  
+uc1     = -5.6e-011     
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.8  nmos
+level = 54
+lmin    = 2.8e-007      
+lmax    = 5e-007        
+wmin    = 1.2e-006      
+wmax    = 1e-005        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.75419347    
+lvth0   = -5.5747725e-008
+wvth0   = -5.7737207e-008
+pvth0   = 1.824977e-014 
+k1      = 0.95060511    
+lk1     = -9.5597554e-008
+wk1     = 1.0355446e-008
+pk1     = -5.177723e-015
+k2      = 0.013945175   
+lk2     = -3.0232209e-008
+wk2     = 1.9443834e-008
+pk2     = -5.4442735e-015
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12424632   
+lvoff   = 6.8691116e-010
+wvoff   = 3.5791497e-008
+pvoff   = -6.8553733e-015
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.046898182   
+lu0     = 1.7050207e-010
+wu0     = -1.6262868e-008
+pu0     = 4.1983839e-015
+ua      = -6.6207759e-010
+lua     = 2.5458994e-016
+wua     = 5.6335718e-017
+pua     = 1.7471409e-022
+ub      = 3.7962141e-018
+lub     = -3.3240512e-025
+wub     = -1.6693412e-024
+pub     = 4.2239319e-032
+uc      = 2.9436835e-010
+luc     = -6.8059408e-017
+wuc     = -1.6002278e-016
+puc     = 3.2259428e-023
+eu      = 1.67          
+vsat    = 85682.645     
+lvsat   = -0.00034132231
+wvsat   = -0.0068127934 
+pvsat   = 3.4063967e-009
+a0      = 0.10362636    
+la0     = -8.0818182e-010
+ags     = 0.2705431     
+lags    = 3.2753448e-008
+wags    = 1.3273025e-007
+pags    = -6.6365124e-014
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.12424077   
+lketa   = 2.9920384e-008
+wketa   = -4.1694295e-009
+pketa   = 2.0847148e-015
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.20476889    
+lpclm   = -9.798626e-009
+wpclm   = 2.8042187e-007
+ppclm   = -5.8632603e-014
+pdiblc1 = 0.39          
+pdiblc2 = 0.003171      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0036363636  
+ldelta  = 3.1818182e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 2.5953123e-006
+lalpha0 = -2.5435614e-013
+walpha0 = 1.1428461e-013
+palpha0 = -5.7142305e-020
+alpha1  = 0             
+beta0   = 21.140586     
+wbeta0  = -5.6473191e-007
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = -0.59809917   
+lnoff   = 1.2990496e-006
+wnoff   = 3.065757e-006 
+pnoff   = -1.5328785e-012
+voffcv  = 0.22872521    
+lvoffcv = -1.118626e-007
+wvoffcv = -2.6399574e-007
+pvoffcv = 1.3199787e-013
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.28115299   
+lkt1    = -1.0099496e-008
+wkt1    = -1.2105482e-007
+pkt1    = 3.5188078e-014
+kt1l    = 0             
+kt2     = -0.025449687  
+lkt2    = 9.6575269e-010
+wkt2    = 8.9970236e-009
+pkt2    = -3.1602845e-015
+ute     = -1.5701136    
+wute    = 2.0073409e-007
+ua1     = 1.675e-009    
+ub1     = -5.3788142e-018
+lub1    = 4.827456e-025 
+wub1    = 2.1072821e-024
+pub1    = -3.1500653e-031
+uc1     = -2.2938539e-010
+luc1    = 4.973267e-017 
+wuc1    = 2.0459475e-016
+puc1    = -5.8684551e-023
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.9  nmos
+level = 54
+lmin    = 5e-007        
+lmax    = 1.2e-006      
+wmin    = 1.2e-006      
+wmax    = 1e-005        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.66260505    
+lvth0   = -9.953513e-009
+wvth0   = 3.6992425e-009
+pvth0   = -1.2468455e-014
+k1      = 0.75941       
+k2      = 0.017155231   
+lk2     = -3.1837237e-008
+wk2     = -6.1109193e-009
+pk2     = 7.3331031e-015
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.10253679   
+lvoff   = -1.0167857e-008
+wvoff   = -1.5771964e-008
+pvoff   = 1.8926357e-014
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.038465008   
+lu0     = 4.387089e-009 
+wu0     = -8.4602728e-009
+pu0     = 2.9708645e-016
+ua      = -9.289245e-010
+lua     = 3.880134e-016 
+wua     = -2.8983135e-016
+pua     = 3.4779762e-022
+ub      = 3.4725304e-018
+lub     = -1.7056325e-025
+wub     = -6.6767982e-025
+pub     = -4.5859137e-031
+uc      = 1.5722431e-010
+luc     = 5.1261039e-019
+wuc     = -8.5272224e-017
+puc     = -5.1158517e-024
+eu      = 1.67          
+vsat    = 85000         
+a0      = 0.57970277    
+la0     = -2.3884638e-007
+wa0     = 4.6802014e-007
+pa0     = -2.3401007e-013
+ags     = 0.63340774    
+lags    = -1.4867887e-007
+wags    = -1.6558842e-007
+pags    = 8.279421e-014 
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.043888571  
+lketa   = -1.0255714e-008
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.047719      
+lpclm   = 6.8726318e-008
+wpclm   = 1.7942187e-007
+ppclm   = -8.1325983e-015
+pdiblc1 = 0.39          
+pdiblc2 = 0.001359      
+lpdiblc2= 9.06e-010     
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0014285714  
+ldelta  = 4.2857143e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 6.7040286e-006
+lalpha0 = -2.3087143e-012
+alpha1  = 0             
+beta0   = 21.043581     
+lbeta0  = 4.8502597e-008
+wbeta0  = 4.0337993e-007
+pbeta0  = -4.8405592e-013
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.30297354   
+lkt1    = 8.1077922e-010
+wkt1    = -9.3348999e-008
+pkt1    = 2.1335166e-014
+kt1l    = 0             
+kt2     = -0.021799026  
+lkt2    = -8.5957792e-010
+wkt2    = -5.9264351e-009
+pkt2    = 4.3014448e-015
+ute     = -1.5701136    
+wute    = 2.0073409e-007
+ua1     = 1.675e-009    
+ub1     = -3.0334126e-018
+lub1    = -6.899552e-025
+wub1    = 3.2333483e-025
+pub1    = 5.7696713e-031
+uc1     = -1.4511739e-010
+luc1    = 7.5986727e-018
+wuc1    = 6.1137104e-017
+puc1    = 1.3044275e-023
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.10  nmos
+level = 54
+lmin    = 1.2e-006      
+lmax    = 1e-005        
+wmin    = 1.2e-006      
+wmax    = 1e-005        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.64815901    
+lvth0   = 7.3817355e-009
+wvth0   = -2.7981116e-009
+pvth0   = -4.6716298e-015
+k1      = 0.79747612    
+lk1     = -4.5679339e-008
+wk1     = -3.0414256e-009
+pk1     = 3.6497107e-015
+k2      = -0.0074231864 
+lk2     = -2.3431364e-009
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12197591   
+lvoff   = 1.3159091e-008
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.040494054   
+lu0     = 1.9522345e-009
+wu0     = -5.9939808e-009
+pu0     = -2.662464e-015
+ua      = -8.1072595e-010
+lua     = 2.4617513e-016
+wua     = 1.9601988e-017
+pua     = -2.3522386e-023
+ub      = 3.1895805e-018
+lub     = 1.6897655e-025
+wub     = -3.2156993e-025
+pub     = -8.7392324e-031
+uc      = 1.0432829e-010
+luc     = 6.3987831e-017
+wuc     = -1.6449976e-017
+puc     = -8.7702549e-023
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.175342      
+la0     = -9.536135e-007
+wa0     = 6.8460666e-008
+pa0     = 2.454613e-013 
+ags     = 0.26729169    
+lags    = 2.9066039e-007
+wags    = 4.3516718e-009
+pags    = -1.211339e-013
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.021025909  
+lketa   = -3.7690909e-008
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.23344442    
+lpclm   = -1.5414418e-007
+wpclm   = -2.3542459e-008
+ppclm   = 2.3542459e-013
+pdiblc1 = 0.39          
+pdiblc2 = 0.00064013636 
+lpdiblc2= 1.7686364e-009
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0027272727  
+ldelta  = 2.7272727e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 9.0929986e-005
+lalpha0 = -1.0337986e-010
+alpha1  = 0             
+beta0   = 24.512311     
+lbeta0  = -4.1139731e-006
+wbeta0  = -3.6192965e-007
+pbeta0  = 4.3431558e-013
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2.128874      
+lnoff   = -1.5464876e-007
+wnoff   = -1.5207128e-007
+pnoff   = 1.8248554e-013
+voffcv  = -0.065880682  
+lvoffcv = 8.5056818e-008
+wvoffcv = 8.3639205e-008
+pvoffcv = -1.0036705e-013
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.31506405   
+lkt1    = 1.5319401e-008
+wkt1    = -3.095198e-008
+pkt1    = -5.3541257e-014
+kt1l    = 0             
+kt2     = -0.016812862  
+lkt2    = -6.8429752e-009
+wkt2    = -5.3833233e-009
+pkt2    = 3.6497107e-015
+ute     = -1.5472572    
+lute    = -2.7427686e-008
+wute    = -2.7372831e-008
+pute    = 2.7372831e-013
+ua1     = 1.6533492e-009
+lua1    = 2.5980992e-017
+wua1    = 2.5547975e-017
+pua1    = -3.065757e-023
+ub1     = -2.1483391e-018
+lub1    = -1.7520434e-024
+wub1    = -1.1332474e-024
+pub1    = 2.3248657e-030
+uc1     = -4.4711114e-011
+luc1    = -1.1288886e-016
+wuc1    = -9.8191818e-018
+puc1    = 9.8191818e-023
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.11  nmos
+level = 54
+lmin    = 1e-005        
+lmax    = 5.0001e-005   
+wmin    = 1.2e-006      
+wmax    = 1e-005        
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.64889718    
+wvth0   = -3.2652745e-009
+k1      = 0.79290818    
+wk1     = -2.6764545e-009
+k2      = -0.0076575    
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12066      
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.040689277   
+wu0     = -6.2602272e-009
+ua      = -7.8610843e-010
+wua     = 1.7249749e-017
+ub      = 3.2064782e-018
+wub     = -4.0896225e-025
+uc      = 1.1072708e-010
+wuc     = -2.5220231e-017
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.0799807     
+wa0     = 9.3006796e-008
+ags     = 0.29635773    
+wags    = -7.7617182e-009
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.024795     
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.21803       
+pdiblc1 = 0.39          
+pdiblc2 = 0.000817      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.003         
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 8.0592e-005   
+alpha1  = 0             
+beta0   = 24.100914     
+wbeta0  = -3.1849809e-007
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2.1134091     
+wnoff   = -1.3382273e-007
+voffcv  = -0.057375     
+wvoffcv = 7.36025e-008  
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.31353211   
+wkt1    = -3.6306106e-008
+kt1l    = 0             
+kt2     = -0.017497159  
+wkt2    = -5.0183523e-009
+ute     = -1.55         
+ua1     = 1.6559473e-009
+wua1    = 2.2482218e-017
+ub1     = -2.3235434e-018
+wub1    = -9.0076078e-025
+uc1     = -5.6e-011     
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.12  nmos
+level = 54
+lmin    = 2.8e-007      
+lmax    = 5e-007        
+wmin    = 1e-005        
+wmax    = 0.000100001   
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 3e-008        
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.74840818    
+lvth0   = -5.3919091e-008
+k1      = 0.95164273    
+lk1     = -9.6116364e-008
+k2      = 0.015893454   
+lk2     = -3.0777727e-008
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12066      
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.045268636   
+lu0     = 5.9118182e-010
+ua      = -6.5643273e-010
+lua     = 2.7209636e-016
+ub      = 3.6289455e-018
+lub     = -3.2817273e-025
+uc      = 2.78334e-010  
+luc     = -6.4827e-017  
+eu      = 1.67          
+vsat    = 85000         
+a0      = 0.13211844    
+la0     = -1.5054221e-008
+wa0     = -2.8435094e-007
+pa0     = 1.4217547e-013
+ags     = 0.46155061    
+lags    = -6.2750307e-008
+wags    = -1.7735247e-006
+pags    = 8.8676235e-013
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.12105603   
+lketa   = 2.8328017e-008
+wketa   = -3.5953066e-008
+pketa   = 1.7976533e-014
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.23286727    
+lpclm   = -1.5673636e-008
+pdiblc1 = 0.39          
+pdiblc2 = 0.003171      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0036363636  
+ldelta  = 3.1818182e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 2.6067636e-006
+lalpha0 = -2.6008182e-013
+alpha1  = 0             
+beta0   = 21.084        
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 2.3e-010      
+cgdo    = 2.3e-010      
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = -0.29090909   
+lnoff   = 1.1454545e-006
+voffcv  = 0.20227273    
+lvoffcv = -9.8636364e-008
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.29328273   
+lkt1    = -6.5736364e-009
+kt1l    = 0             
+kt2     = -0.024548182  
+lkt2    = 6.4909091e-010
+ute     = -1.55         
+ua1     = 1.675e-009    
+ub1     = -5.1676636e-018
+lub1    = 4.5118182e-025
+uc1     = -2.0888491e-010
+luc1    = 4.3852454e-017
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.13  nmos
+level = 54
+lmin    = 5e-007        
+lmax    = 1.2e-006      
+wmin    = 1e-005        
+wmax    = 0.000100001   
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.66297571    
+lvth0   = -1.1202857e-008
+k1      = 0.75941       
+k2      = 0.016542914   
+lk2     = -3.1102457e-008
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.10411714   
+lvoff   = -8.2714286e-009
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.037617286   
+lu0     = 4.4168571e-009
+ua      = -9.5796571e-010
+lua     = 4.2286286e-016
+ub      = 3.4056286e-018
+lub     = -2.1651429e-025
+uc      = 1.4868e-010   
+eu      = 1.67          
+vsat    = 85000         
+a0      = 0.62659857    
+la0     = -2.6229429e-007
+ags     = 0.61681571    
+lags    = -1.4038286e-007
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.043888571  
+lketa   = -1.0255714e-008
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.065697143   
+lpclm   = 6.7911429e-008
+pdiblc1 = 0.39          
+pdiblc2 = 0.001359      
+lpdiblc2= 9.06e-010     
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0014285714  
+ldelta  = 4.2857143e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 6.7040286e-006
+lalpha0 = -2.3087143e-012
+alpha1  = 0             
+beta0   = 21.084        
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2             
+voffcv  = 0.005         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.31232714   
+lkt1    = 2.9485714e-009
+kt1l    = 0             
+kt2     = -0.022392857  
+lkt2    = -4.2857143e-010
+ute     = -1.55         
+ua1     = 1.675e-009    
+ub1     = -3.0010143e-018
+lub1    = -6.3214286e-025
+uc1     = -1.3899143e-010
+luc1    = 8.9057143e-018
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.14  nmos
+level = 54
+lmin    = 1.2e-006      
+lmax    = 1e-005        
+wmin    = 1e-005        
+wmax    = 0.000100001   
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 0             
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.64787864    
+lvth0   = 6.9136364e-009
+k1      = 0.79717136    
+lk1     = -4.5313636e-008
+k2      = -0.0074231864 
+lk2     = -2.3431364e-009
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12197591   
+lvoff   = 1.3159091e-008
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.039893455   
+lu0     = 1.6854546e-009
+ua      = -8.0876182e-010
+lua     = 2.4381818e-016
+ub      = 3.1573591e-018
+lub     = 8.1409091e-026
+uc      = 1.0268e-010   
+luc     = 5.52e-017     
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.1822018     
+la0     = -9.2901818e-007
+ags     = 0.26772773    
+lags    = 2.7852273e-007
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.021025909  
+lketa   = -3.7690909e-008
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.23108545    
+lpclm   = -1.3055455e-007
+pdiblc1 = 0.39          
+pdiblc2 = 0.00064013636 
+lpdiblc2= 1.7686364e-009
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.0027272727  
+ldelta  = 2.7272727e-009
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 9.0929986e-005
+lalpha0 = -1.0337986e-010
+alpha1  = 0             
+beta0   = 24.476046     
+lbeta0  = -4.0704545e-006
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 1e-010        
+cgdo    = 1e-010        
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2.1136364     
+lnoff   = -1.3636364e-007
+voffcv  = -0.0575       
+lvoffcv = 7.5e-008      
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.31816545   
+lkt1    = 9.9545454e-009
+kt1l    = 0             
+kt2     = -0.017352273  
+lkt2    = -6.4772727e-009
+ute     = -1.55         
+ua1     = 1.6559091e-009
+lua1    = 2.2909091e-017
+ub1     = -2.2618909e-018
+lub1    = -1.5190909e-024
+uc1     = -4.5695e-011  
+luc1    = -1.0305e-016  
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.model  nmos_3p3.15  nmos
+level = 54
+lmin    = 1e-005        
+lmax    = 5.0001e-005   
+wmin    = 1e-005        
+wmax    = 0.000100001   
+version = 4.5           
+binunit = 2             
+paramchk= 1             
+mobmod  = 0             
+capmod  = 2             
+igcmod  = 0             
+igbmod  = 0             
+geomod  = 0             
+diomod  = 1             
+rdsmod  = 0             
+rbodymod= 0             
+rgatemod= 0             
+permod  = 1             
+acnqsmod= 0             
+trnqsmod= 0             
+tnom    = 25            
+toxe    = 8e-009        
+toxp    = 8e-009        
+toxm    = 8e-009        
+epsrox  = 3.9           
+wint    = 1e-008        
+lint    = 0             
+ll      = 0             
+wl      = 0             
+lln     = 1             
+wln     = 1             
+lw      = 0             
+ww      = 0             
+lwn     = 1             
+wwn     = 1             
+lwl     = 0             
+wwl     = 0             
+xl      = 0             
+xw      = 0             
+dlc     = 3e-008        
+dwc     = 0             
+xpart   = 0             
+toxref  = 8e-009        
+dlcig   = 1.5e-007      
+vth0    = 0.64857       
+k1      = 0.79264       
+k2      = -0.0076575    
+k3      = 0             
+k3b     = 0             
+w0      = 5e-007        
+dvt0    = 0             
+dvt1    = 0.53          
+dvt2    = 0             
+dvt0w   = 0             
+dvt1w   = 0             
+dvt2w   = 0             
+dsub    = 0.5           
+minv    = -0.25         
+voffl   = 0             
+dvtp0   = 0             
+dvtp1   = 0             
+lpe0    = 1.1e-007      
+lpeb    = 0             
+vbm     = -3            
+xj      = 1e-007        
+ngate   = 6e+019        
+ndep    = 3e+017        
+nsd     = 1e+020        
+phin    = 0.07          
+cdsc    = 0             
+cdscb   = 0             
+cdscd   = 0             
+cit     = 0             
+voff    = -0.12066      
+nfactor = 1             
+eta0    = 0.75          
+etab    = -0.32         
+u0      = 0.040062      
+ua      = -7.8438e-010  
+ub      = 3.1655e-018   
+uc      = 1.082e-010    
+eu      = 1.67          
+vsat    = 85000         
+a0      = 1.0893        
+ags     = 0.29558       
+a1      = 0             
+a2      = 1             
+b0      = 0             
+b1      = 0             
+keta    = -0.024795     
+dwg     = 0             
+dwb     = 0             
+pclm    = 0.21803       
+pdiblc1 = 0.39          
+pdiblc2 = 0.000817      
+pdiblcb = 0.2           
+drout   = 0.56          
+pvag    = 0             
+delta   = 0.003         
+pscbe1  = 6.6469e+008   
+pscbe2  = 1.638e-005    
+fprout  = 0             
+pdits   = 0             
+pditsd  = 0             
+pditsl  = 0             
+rsh     = 7             
+rdsw    = 530           
+rdswmin = 50            
+rdwmin  = 0             
+rswmin  = 0             
+prwg    = 0             
+prwb    = 0             
+wr      = 1             
+alpha0  = 8.0592e-005   
+alpha1  = 0             
+beta0   = 24.069        
+agidl   = 1.3268e-010   
+bgidl   = 1.8961e+009   
+cgidl   = 0.5           
+egidl   = 0.8           
+cgso    = 2.3e-010      
+cgdo    = 2.3e-010      
+cgbo    = 1e-013        
+cgdl    = 1e-010        
+cgsl    = 1e-010        
+clc     = 1e-007        
+cle     = 0.6           
+cf      = 0             
+ckappas = 0.6           
+ckappad = 0.6           
+vfbcv   = -1            
+acde    = 0.6           
+moin    = 15            
+noff    = 2.1           
+voffcv  = -0.05         
+tvoff   = 0.001         
+ltvoff  = 0             
+wtvoff  = 0             
+ptvoff  = 0             
+kt1     = -0.31717      
+kt1l    = 0             
+kt2     = -0.018        
+ute     = -1.55         
+ua1     = 1.6582e-009   
+ub1     = -2.4138e-018  
+uc1     = -5.6e-011     
+prt     = 0             
+at      = 23000         
+fnoimod = 1             
+tnoimod = 0             
+em      = 4.1e+007      
+ef      = 0.95          
+noia    = nmos_3p3_noia  
+noib    = nmos_3p3_noib  
+noic    = nmos_3p3_noic  
+ntnoi   = 1             
+jss     = 2.2959e-007   
+jsws    = 2.1207e-013   
+jswgs   = 0             
+njs     = 1.01          
+ijthsfwd= 0.1           
+ijthsrev= 0.1           
+pbs     = 0.70172       
+cjs     = 0.00096797    
+mjs     = 0.32071       
+pbsws   = 0.8062        
+cjsws   = 1.5663e-010   
+mjsws   = 0.1           
+pbswgs  = 0.74743       
+cjswgs  = 5.9903e-010   
+mjswgs  = 0.32059       
+tpb     = 0.0018129     
+tcj     = 0.0009438     
+tpbsw   = 5e-005        
+tcjsw   = 0.00060474    
+tpbswg  = 0.0016872     
+tcjswg  = 0.001         
+xtis    = 3             
+dmcg    = 1.5e-007      
+saref   = 4.4e-007      
+sbref   = 4.4e-007      
+kvth0   = 0             
+ku0     = 0             
+kvsat   = 0             
.title KiCad schematic
V1 Net-_V1-E1_ 0 1
R1 Net-_V1-E1_ out 1k
R2 out 0 2k
.end

* This first line is a comment.
.param mega=1MEG milli=1M one='mega*milli'

.tran 0.1 1
.tran 0.1 1 uic
.tran 0.1 1 0
.tran 0.1 1 0 uic
.tran 0.1 1 0 0.2
.tran 0.1 1 0 0.2 uic

* Title
*.GLOBAL VDD
*.GLOBAL VSS
.OPTION gmin=1e-15
VVDD VDD 0 5.0
VVSS VSS 0 0.0
.INCLUDE "gf180mcu_fd_sc_mcu7t5v0__dffnq_4.ngspice"
CQ Q_tmp 0 1.7205e-13
VQ Q Q_tmp 0
VNW VNW VDD 0
VPW VPW VSS 0

VCLKN CLKN 0 PWL(
+ 000000.0e-12 5.0
+ 050000.0e-12 5.0
+ 051020.0e-12 0.0
+ 100000.0e-12 0.0
+ 101020.0e-12 5.0
+ 400000.0e-12 5.0
+ 401020.0e-12 0.0
+ 500000.0e-12 0.0
+ 501020.0e-12 5.0
+ 600000.0e-12 5.0
+ 601020.0e-12 0.0
+ 700000.0e-12 0.0
+ )
VD D 0 PWL(
+ 000000.0e-12 0.0
+ 200000.0e-12 0.0
+ 201020.0e-12 5.0
+ 300000.0e-12 5.0
+ 301020.0e-12 0.0
+ 400000.0e-12 0.0
+ 401020.0e-12 5.0
+ 600000.0e-12 5.0
+ )
.LIB "jlpkg://GF180MCUPDK/sm141064.ngspice" statistical
.TRAN 3.3333333333333e-10 6.0e-7
.END
